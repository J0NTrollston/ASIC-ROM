** sch_path: /home/ttuser/Documents/ASIC-ROM/xschem/testbench.sch
**.subckt testbench
x1 VDD VSS x0 x1 en PC b2 b1 b0 b3 NOR_ROM_2bit
V1 VDD GND 1.8
V2 VSS GND 0
V4 x1 GND 0
V3 x0 GND 1.8
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/ttuser/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /home/ttuser/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice





Ven en 0 PWL (0ms 0V 20ms 0V 22ms 1.8V)
VPC PC 0 PWL(0ms 0V .9ms 0V 1ms 1.8V)
* Ven en 0 PWL (0ms 0V 3ms 0V 3.1ms 1.8V 9.8ms 1.8V 9.9ms 0V )
* VPC PC 0 PWL(0ms 0V .9ms 0V 1ms 1.8V 10ms 1.8V 10.1ms 0V 10.9ms 0V 11ms 1.8V 20ms 1.8V 20.1ms 0V 20.9ms 0V 21ms 1.8V 30ms 1.8V 30.1ms 0V 30.9ms 0V 31ms 1.8V)
* Vx0 x0 0 PWL(0ms 0V 9.9ms 0V 10ms 1.8V 19.9ms 1.8V 20ms 0V 29.9ms 0V 30ms 1.8V )
* Vx1 x1 0 PWL(0ms 0V 9.9ms 0V 10ms 0V 19.9ms 0V 20ms 1.8V)

.control
tran 1us 50ms
write testbench.raw
.endc



**** end user architecture code
**.ends

* expanding   symbol:  NOR_ROM_2bit.sym # of pins=10
** sym_path: /home/ttuser/Documents/ASIC-ROM/xschem/NOR_ROM_2bit.sym
** sch_path: /home/ttuser/Documents/ASIC-ROM/xschem/NOR_ROM_2bit.sch
.subckt NOR_ROM_2bit VDD VSS x0 x1 en PC b1 b2 b0 b3
*.iopin VDD
*.iopin VSS
*.ipin x0
*.opin b3
*.ipin x1
*.opin b2
*.opin b1
*.opin b0
*.ipin PC
*.ipin en
XM4 b0_n D VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 b1_n C VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 b0_n C VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 b2_n B VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 b1_n B VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 b0_n B VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 b0_n A VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 b1_n A VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM13 b2_n A VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM14 b3_n A VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x1 b3_n VGND VNB VPB VPWR b3 sky130_fd_sc_hd__inv_1
x2 b2_n VGND VNB VPB VPWR b2 sky130_fd_sc_hd__inv_1
x3 b1_n VGND VNB VPB VPWR b1 sky130_fd_sc_hd__inv_1
x4 b0_n VGND VNB VPB VPWR b0 sky130_fd_sc_hd__inv_1
x9 x1 VGND VNB VPB VPWR x1_n sky130_fd_sc_hd__inv_1
x10 x0 VGND VNB VPB VPWR x0_n sky130_fd_sc_hd__inv_1
XM1 b3_n PC VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 b2_n PC VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 b1_n PC VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 b0_n PC VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x11 x0_n x1_n en VGND VNB VPB VPWR D sky130_fd_sc_hd__and3_1
x5 x0 x1_n en VGND VNB VPB VPWR C sky130_fd_sc_hd__and3_1
x6 x0_n x1 en VGND VNB VPB VPWR B sky130_fd_sc_hd__and3_1
x7 x0 x1 en VGND VNB VPB VPWR A sky130_fd_sc_hd__and3_1
.ends

.GLOBAL GND
.end
